module mainProcessor();


endmodule