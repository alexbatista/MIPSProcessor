module alu
#(parameter WIDTH=32)
(input [WIDTH-1:0] a, input [WIDTH-1:0]b, input [2:0] sel);


endmodule